magic
tech sky130A
timestamp 1766605324
<< nwell >>
rect -835 1090 -610 1265
rect -475 1015 210 1190
rect 340 955 565 1115
rect 745 1095 970 1270
rect 1105 1020 1790 1195
rect 1920 960 2145 1120
rect 370 940 565 955
rect 1950 945 2145 960
rect 2280 900 2655 1060
rect 790 855 980 860
rect -790 850 -600 855
rect -790 680 -565 850
rect 90 540 530 715
rect 790 685 1015 855
rect 1670 545 2110 720
<< nmos >>
rect -705 955 -690 1055
rect -660 545 -645 645
rect -345 785 -330 885
rect -240 785 -225 885
rect -35 785 -20 885
rect 70 785 85 885
rect 875 960 890 1060
rect 470 805 485 905
rect 920 550 935 650
rect 1235 790 1250 890
rect 1340 790 1355 890
rect 1545 790 1560 890
rect 1650 790 1665 890
rect 2050 810 2065 910
rect 2405 750 2420 850
rect 2510 750 2525 850
rect 210 375 225 475
rect 315 375 330 475
rect 1790 320 1805 420
rect 1895 320 1910 420
<< pmos >>
rect -705 1125 -690 1225
rect -345 1050 -330 1150
rect -240 1050 -225 1150
rect -35 1050 -20 1150
rect 70 1050 85 1150
rect -660 715 -645 815
rect 875 1130 890 1230
rect 470 975 485 1075
rect 1235 1055 1250 1155
rect 1340 1055 1355 1155
rect 1545 1055 1560 1155
rect 1650 1055 1665 1155
rect 920 720 935 820
rect 210 575 225 675
rect 315 575 330 675
rect 2050 980 2065 1080
rect 2405 925 2420 1025
rect 2510 925 2525 1025
rect 1790 580 1805 680
rect 1895 580 1910 680
<< ndiff >>
rect -750 1040 -705 1055
rect -750 970 -740 1040
rect -720 970 -705 1040
rect -750 955 -705 970
rect -690 1040 -645 1055
rect -690 970 -675 1040
rect -655 970 -645 1040
rect -690 955 -645 970
rect -705 630 -660 645
rect -705 560 -695 630
rect -675 560 -660 630
rect -705 545 -660 560
rect -645 630 -600 645
rect -645 560 -630 630
rect -610 560 -600 630
rect -410 870 -345 885
rect -410 800 -380 870
rect -360 800 -345 870
rect -410 785 -345 800
rect -330 870 -240 885
rect -330 800 -315 870
rect -295 800 -275 870
rect -255 800 -240 870
rect -330 785 -240 800
rect -225 870 -180 885
rect -100 870 -35 885
rect -225 800 -210 870
rect -190 800 -180 870
rect -100 800 -70 870
rect -50 800 -35 870
rect -225 785 -180 800
rect -100 785 -35 800
rect -20 870 70 885
rect -20 800 -5 870
rect 15 800 35 870
rect 55 800 70 870
rect -20 785 70 800
rect 85 870 130 885
rect 85 800 100 870
rect 120 800 130 870
rect 830 1045 875 1060
rect 830 975 840 1045
rect 860 975 875 1045
rect 830 960 875 975
rect 890 1045 935 1060
rect 890 975 905 1045
rect 925 975 935 1045
rect 890 960 935 975
rect 425 890 470 905
rect 85 785 130 800
rect 425 820 435 890
rect 455 820 470 890
rect 425 805 470 820
rect 485 890 530 905
rect 485 820 500 890
rect 520 820 530 890
rect 485 805 530 820
rect 875 635 920 650
rect -645 545 -600 560
rect 875 565 885 635
rect 905 565 920 635
rect 875 550 920 565
rect 935 635 980 650
rect 935 565 950 635
rect 970 565 980 635
rect 1170 875 1235 890
rect 1170 805 1200 875
rect 1220 805 1235 875
rect 1170 790 1235 805
rect 1250 875 1340 890
rect 1250 805 1265 875
rect 1285 805 1305 875
rect 1325 805 1340 875
rect 1250 790 1340 805
rect 1355 875 1400 890
rect 1480 875 1545 890
rect 1355 805 1370 875
rect 1390 805 1400 875
rect 1480 805 1510 875
rect 1530 805 1545 875
rect 1355 790 1400 805
rect 1480 790 1545 805
rect 1560 875 1650 890
rect 1560 805 1575 875
rect 1595 805 1615 875
rect 1635 805 1650 875
rect 1560 790 1650 805
rect 1665 875 1710 890
rect 1665 805 1680 875
rect 1700 805 1710 875
rect 2005 895 2050 910
rect 1665 790 1710 805
rect 2005 825 2015 895
rect 2035 825 2050 895
rect 2005 810 2050 825
rect 2065 895 2110 910
rect 2065 825 2080 895
rect 2100 825 2110 895
rect 2065 810 2110 825
rect 2360 835 2405 850
rect 2360 765 2370 835
rect 2390 765 2405 835
rect 2360 750 2405 765
rect 2420 835 2510 850
rect 2420 765 2435 835
rect 2455 765 2475 835
rect 2495 765 2510 835
rect 2420 750 2510 765
rect 2525 835 2570 850
rect 2525 765 2540 835
rect 2560 765 2570 835
rect 2525 750 2570 765
rect 935 550 980 565
rect 145 460 210 475
rect 145 390 175 460
rect 195 390 210 460
rect 145 375 210 390
rect 225 460 315 475
rect 225 390 240 460
rect 260 390 280 460
rect 300 390 315 460
rect 225 375 315 390
rect 330 460 375 475
rect 330 390 345 460
rect 365 390 375 460
rect 330 375 375 390
rect 1725 405 1790 420
rect 1725 335 1755 405
rect 1775 335 1790 405
rect 1725 320 1790 335
rect 1805 405 1895 420
rect 1805 335 1820 405
rect 1840 335 1860 405
rect 1880 335 1895 405
rect 1805 320 1895 335
rect 1910 405 1955 420
rect 1910 335 1925 405
rect 1945 335 1955 405
rect 1910 320 1955 335
<< pdiff >>
rect -750 1210 -705 1225
rect -750 1140 -740 1210
rect -720 1140 -705 1210
rect -750 1125 -705 1140
rect -690 1210 -645 1225
rect -690 1140 -675 1210
rect -655 1140 -645 1210
rect 830 1215 875 1230
rect -690 1125 -645 1140
rect -390 1135 -345 1150
rect -390 1065 -380 1135
rect -360 1065 -345 1135
rect -390 1050 -345 1065
rect -330 1135 -240 1150
rect -330 1065 -315 1135
rect -295 1065 -275 1135
rect -255 1065 -240 1135
rect -330 1050 -240 1065
rect -225 1135 -180 1150
rect -95 1135 -35 1150
rect -225 1065 -210 1135
rect -190 1065 -180 1135
rect -95 1065 -70 1135
rect -50 1065 -35 1135
rect -225 1050 -180 1065
rect -95 1050 -35 1065
rect -20 1135 70 1150
rect -20 1065 -5 1135
rect 15 1065 35 1135
rect 55 1065 70 1135
rect -20 1050 70 1065
rect 85 1135 150 1150
rect 85 1065 100 1135
rect 120 1065 150 1135
rect 85 1050 150 1065
rect -705 800 -660 815
rect -705 730 -695 800
rect -675 730 -660 800
rect -705 715 -660 730
rect -645 800 -600 815
rect -645 730 -630 800
rect -610 730 -600 800
rect -645 715 -600 730
rect 830 1145 840 1215
rect 860 1145 875 1215
rect 830 1130 875 1145
rect 890 1215 935 1230
rect 890 1145 905 1215
rect 925 1145 935 1215
rect 890 1130 935 1145
rect 1190 1140 1235 1155
rect 425 1060 470 1075
rect 425 990 435 1060
rect 455 990 470 1060
rect 425 975 470 990
rect 485 1060 530 1075
rect 485 990 500 1060
rect 520 990 530 1060
rect 485 975 530 990
rect 1190 1070 1200 1140
rect 1220 1070 1235 1140
rect 1190 1055 1235 1070
rect 1250 1140 1340 1155
rect 1250 1070 1265 1140
rect 1285 1070 1305 1140
rect 1325 1070 1340 1140
rect 1250 1055 1340 1070
rect 1355 1140 1400 1155
rect 1485 1140 1545 1155
rect 1355 1070 1370 1140
rect 1390 1070 1400 1140
rect 1485 1070 1510 1140
rect 1530 1070 1545 1140
rect 1355 1055 1400 1070
rect 1485 1055 1545 1070
rect 1560 1140 1650 1155
rect 1560 1070 1575 1140
rect 1595 1070 1615 1140
rect 1635 1070 1650 1140
rect 1560 1055 1650 1070
rect 1665 1140 1730 1155
rect 1665 1070 1680 1140
rect 1700 1070 1730 1140
rect 1665 1055 1730 1070
rect 875 805 920 820
rect 875 735 885 805
rect 905 735 920 805
rect 875 720 920 735
rect 935 805 980 820
rect 935 735 950 805
rect 970 735 980 805
rect 935 720 980 735
rect 165 660 210 675
rect 165 590 175 660
rect 195 590 210 660
rect 165 575 210 590
rect 225 660 315 675
rect 225 590 240 660
rect 260 590 280 660
rect 300 590 315 660
rect 225 575 315 590
rect 330 660 375 675
rect 330 590 345 660
rect 365 590 375 660
rect 330 575 375 590
rect 2005 1065 2050 1080
rect 2005 995 2015 1065
rect 2035 995 2050 1065
rect 2005 980 2050 995
rect 2065 1065 2110 1080
rect 2065 995 2080 1065
rect 2100 995 2110 1065
rect 2065 980 2110 995
rect 2360 1010 2405 1025
rect 2360 940 2370 1010
rect 2390 940 2405 1010
rect 2360 925 2405 940
rect 2420 1010 2510 1025
rect 2420 940 2435 1010
rect 2455 940 2475 1010
rect 2495 940 2510 1010
rect 2420 925 2510 940
rect 2525 1010 2590 1025
rect 2525 940 2540 1010
rect 2560 940 2590 1010
rect 2525 925 2590 940
rect 1745 665 1790 680
rect 1745 595 1755 665
rect 1775 595 1790 665
rect 1745 580 1790 595
rect 1805 665 1895 680
rect 1805 595 1820 665
rect 1840 595 1860 665
rect 1880 595 1895 665
rect 1805 580 1895 595
rect 1910 665 1955 680
rect 1910 595 1925 665
rect 1945 595 1955 665
rect 1910 580 1955 595
<< ndiffc >>
rect -740 970 -720 1040
rect -675 970 -655 1040
rect -695 560 -675 630
rect -630 560 -610 630
rect -380 800 -360 870
rect -315 800 -295 870
rect -275 800 -255 870
rect -210 800 -190 870
rect -70 800 -50 870
rect -5 800 15 870
rect 35 800 55 870
rect 100 800 120 870
rect 840 975 860 1045
rect 905 975 925 1045
rect 435 820 455 890
rect 500 820 520 890
rect 885 565 905 635
rect 950 565 970 635
rect 1200 805 1220 875
rect 1265 805 1285 875
rect 1305 805 1325 875
rect 1370 805 1390 875
rect 1510 805 1530 875
rect 1575 805 1595 875
rect 1615 805 1635 875
rect 1680 805 1700 875
rect 2015 825 2035 895
rect 2080 825 2100 895
rect 2370 765 2390 835
rect 2435 765 2455 835
rect 2475 765 2495 835
rect 2540 765 2560 835
rect 175 390 195 460
rect 240 390 260 460
rect 280 390 300 460
rect 345 390 365 460
rect 1755 335 1775 405
rect 1820 335 1840 405
rect 1860 335 1880 405
rect 1925 335 1945 405
<< pdiffc >>
rect -740 1140 -720 1210
rect -675 1140 -655 1210
rect -380 1065 -360 1135
rect -315 1065 -295 1135
rect -275 1065 -255 1135
rect -210 1065 -190 1135
rect -70 1065 -50 1135
rect -5 1065 15 1135
rect 35 1065 55 1135
rect 100 1065 120 1135
rect -695 730 -675 800
rect -630 730 -610 800
rect 840 1145 860 1215
rect 905 1145 925 1215
rect 435 990 455 1060
rect 500 990 520 1060
rect 1200 1070 1220 1140
rect 1265 1070 1285 1140
rect 1305 1070 1325 1140
rect 1370 1070 1390 1140
rect 1510 1070 1530 1140
rect 1575 1070 1595 1140
rect 1615 1070 1635 1140
rect 1680 1070 1700 1140
rect 885 735 905 805
rect 950 735 970 805
rect 175 590 195 660
rect 240 590 260 660
rect 280 590 300 660
rect 345 590 365 660
rect 2015 995 2035 1065
rect 2080 995 2100 1065
rect 2370 940 2390 1010
rect 2435 940 2455 1010
rect 2475 940 2495 1010
rect 2540 940 2560 1010
rect 1755 595 1775 665
rect 1820 595 1840 665
rect 1860 595 1880 665
rect 1925 595 1945 665
<< psubdiff >>
rect -790 1040 -750 1055
rect -790 970 -780 1040
rect -760 970 -750 1040
rect -790 955 -750 970
rect -745 630 -705 645
rect -745 560 -735 630
rect -715 560 -705 630
rect -745 545 -705 560
rect -450 870 -410 885
rect -450 800 -440 870
rect -420 800 -410 870
rect -450 785 -410 800
rect -180 870 -100 885
rect -180 800 -170 870
rect -150 800 -130 870
rect -110 800 -100 870
rect -180 785 -100 800
rect 130 870 170 885
rect 130 800 140 870
rect 160 800 170 870
rect 790 1045 830 1060
rect 790 975 800 1045
rect 820 975 830 1045
rect 790 960 830 975
rect 385 890 425 905
rect 130 785 170 800
rect 385 820 395 890
rect 415 820 425 890
rect 385 805 425 820
rect 835 635 875 650
rect 835 565 845 635
rect 865 565 875 635
rect 835 550 875 565
rect 1130 875 1170 890
rect 1130 805 1140 875
rect 1160 805 1170 875
rect 1130 790 1170 805
rect 1400 875 1480 890
rect 1400 805 1410 875
rect 1430 805 1450 875
rect 1470 805 1480 875
rect 1400 790 1480 805
rect 1710 875 1750 890
rect 1710 805 1720 875
rect 1740 805 1750 875
rect 1965 895 2005 910
rect 1710 790 1750 805
rect 1965 825 1975 895
rect 1995 825 2005 895
rect 1965 810 2005 825
rect 2320 835 2360 850
rect 2320 765 2330 835
rect 2350 765 2360 835
rect 2320 750 2360 765
rect 2570 835 2610 850
rect 2570 765 2580 835
rect 2600 765 2610 835
rect 2570 750 2610 765
rect 105 460 145 475
rect 105 390 115 460
rect 135 390 145 460
rect 105 375 145 390
rect 375 460 415 475
rect 375 390 385 460
rect 405 390 415 460
rect 375 375 415 390
rect 1685 405 1725 420
rect 1685 335 1695 405
rect 1715 335 1725 405
rect 1685 320 1725 335
rect 1955 405 1995 420
rect 1955 335 1965 405
rect 1985 335 1995 405
rect 1955 320 1995 335
<< nsubdiff >>
rect -790 1210 -750 1225
rect -790 1140 -780 1210
rect -760 1140 -750 1210
rect -790 1125 -750 1140
rect 790 1215 830 1230
rect -430 1135 -390 1150
rect -430 1065 -420 1135
rect -400 1065 -390 1135
rect -430 1050 -390 1065
rect -180 1135 -95 1150
rect -180 1065 -170 1135
rect -150 1065 -130 1135
rect -110 1065 -95 1135
rect -180 1050 -95 1065
rect 150 1135 190 1150
rect 150 1065 160 1135
rect 180 1065 190 1135
rect 150 1050 190 1065
rect -745 800 -705 815
rect -745 730 -735 800
rect -715 730 -705 800
rect -745 715 -705 730
rect 790 1145 800 1215
rect 820 1145 830 1215
rect 790 1130 830 1145
rect 1150 1140 1190 1155
rect 385 1060 425 1075
rect 385 990 395 1060
rect 415 990 425 1060
rect 385 975 425 990
rect 1150 1070 1160 1140
rect 1180 1070 1190 1140
rect 1150 1055 1190 1070
rect 1400 1140 1485 1155
rect 1400 1070 1410 1140
rect 1430 1070 1450 1140
rect 1470 1070 1485 1140
rect 1400 1055 1485 1070
rect 1730 1140 1770 1155
rect 1730 1070 1740 1140
rect 1760 1070 1770 1140
rect 1730 1055 1770 1070
rect 835 805 875 820
rect 835 735 845 805
rect 865 735 875 805
rect 835 720 875 735
rect 125 660 165 675
rect 125 590 135 660
rect 155 590 165 660
rect 125 575 165 590
rect 375 660 415 675
rect 375 590 385 660
rect 405 590 415 660
rect 375 575 415 590
rect 1965 1065 2005 1080
rect 1965 995 1975 1065
rect 1995 995 2005 1065
rect 1965 980 2005 995
rect 2320 1010 2360 1025
rect 2320 940 2330 1010
rect 2350 940 2360 1010
rect 2320 925 2360 940
rect 2590 1010 2630 1025
rect 2590 940 2600 1010
rect 2620 940 2630 1010
rect 2590 925 2630 940
rect 1705 665 1745 680
rect 1705 595 1715 665
rect 1735 595 1745 665
rect 1705 580 1745 595
rect 1955 665 1995 680
rect 1955 595 1965 665
rect 1985 595 1995 665
rect 1955 580 1995 595
<< psubdiffcont >>
rect -780 970 -760 1040
rect -735 560 -715 630
rect -440 800 -420 870
rect -170 800 -150 870
rect -130 800 -110 870
rect 140 800 160 870
rect 800 975 820 1045
rect 395 820 415 890
rect 845 565 865 635
rect 1140 805 1160 875
rect 1410 805 1430 875
rect 1450 805 1470 875
rect 1720 805 1740 875
rect 1975 825 1995 895
rect 2330 765 2350 835
rect 2580 765 2600 835
rect 115 390 135 460
rect 385 390 405 460
rect 1695 335 1715 405
rect 1965 335 1985 405
<< nsubdiffcont >>
rect -780 1140 -760 1210
rect -420 1065 -400 1135
rect -170 1065 -150 1135
rect -130 1065 -110 1135
rect 160 1065 180 1135
rect -735 730 -715 800
rect 800 1145 820 1215
rect 395 990 415 1060
rect 1160 1070 1180 1140
rect 1410 1070 1430 1140
rect 1450 1070 1470 1140
rect 1740 1070 1760 1140
rect 845 735 865 805
rect 135 590 155 660
rect 385 590 405 660
rect 1975 995 1995 1065
rect 2330 940 2350 1010
rect 2600 940 2620 1010
rect 1715 595 1735 665
rect 1965 595 1985 665
<< poly >>
rect -705 1225 -690 1240
rect 875 1230 890 1245
rect -345 1190 285 1205
rect -345 1150 -330 1190
rect -240 1150 -225 1165
rect -35 1150 -20 1165
rect 70 1150 85 1165
rect -705 1080 -690 1125
rect -835 1065 -690 1080
rect -835 1045 -800 1065
rect -705 1055 -690 1065
rect -705 940 -690 955
rect -705 925 -480 940
rect -550 865 -520 875
rect -550 845 -545 865
rect -525 845 -520 865
rect -550 835 -520 845
rect -660 815 -645 830
rect -660 670 -645 715
rect -790 655 -645 670
rect -790 635 -755 655
rect -660 645 -645 655
rect -540 615 -525 835
rect -495 735 -480 925
rect -345 885 -330 1050
rect -240 885 -225 1050
rect -35 885 -20 1050
rect 70 885 85 1050
rect 270 880 285 1190
rect 1235 1195 1865 1210
rect 1235 1155 1250 1195
rect 1340 1155 1355 1170
rect 1545 1155 1560 1170
rect 1650 1155 1665 1170
rect 470 1075 485 1090
rect 875 1085 890 1130
rect 645 1070 890 1085
rect 315 935 355 945
rect 470 935 485 975
rect 645 945 665 1070
rect 875 1060 890 1070
rect 875 945 890 960
rect 315 915 325 935
rect 345 915 485 935
rect 315 905 355 915
rect 470 905 485 915
rect 635 935 675 945
rect 635 915 645 935
rect 665 915 675 935
rect 875 930 1100 945
rect 635 905 675 915
rect 270 865 330 880
rect -345 735 -330 785
rect -495 720 -330 735
rect -355 675 -325 685
rect -240 675 -225 785
rect -35 725 -20 785
rect -355 655 -350 675
rect -330 655 -225 675
rect -200 710 -20 725
rect -355 645 -325 655
rect -200 615 -185 710
rect 70 685 85 785
rect -540 600 -185 615
rect -145 670 85 685
rect 210 675 225 690
rect 315 675 330 865
rect 1030 870 1060 880
rect 1030 850 1035 870
rect 1055 850 1060 870
rect 1030 840 1060 850
rect 920 820 935 835
rect 470 790 485 805
rect 640 675 675 685
rect 920 675 935 720
rect -145 575 -130 670
rect 640 660 935 675
rect 640 650 675 660
rect 920 650 935 660
rect -540 560 -130 575
rect -660 520 -645 545
rect -540 520 -525 560
rect -145 540 -130 560
rect 210 540 225 575
rect -145 525 225 540
rect -660 505 -525 520
rect 210 475 225 525
rect 315 475 330 575
rect 1040 620 1055 840
rect 1085 740 1100 930
rect 1235 890 1250 1055
rect 1340 890 1355 1055
rect 1545 890 1560 1055
rect 1650 890 1665 1055
rect 1850 885 1865 1195
rect 2050 1080 2065 1095
rect 2405 1025 2420 1040
rect 2510 1025 2525 1040
rect 1895 940 1935 950
rect 2050 940 2065 980
rect 1895 920 1905 940
rect 1925 920 2065 940
rect 1895 910 1935 920
rect 2050 910 2065 920
rect 1850 870 1910 885
rect 1235 740 1250 790
rect 1085 725 1250 740
rect 1225 680 1255 690
rect 1340 680 1355 790
rect 1545 730 1560 790
rect 1225 660 1230 680
rect 1250 660 1355 680
rect 1380 715 1560 730
rect 1225 650 1255 660
rect 1380 620 1395 715
rect 1650 690 1665 790
rect 1040 605 1395 620
rect 1435 675 1665 690
rect 1790 680 1805 695
rect 1895 680 1910 870
rect 2405 850 2420 925
rect 2510 850 2525 925
rect 2050 795 2065 810
rect 1435 580 1450 675
rect 2405 675 2420 750
rect 2400 665 2430 675
rect 2510 665 2525 750
rect 2400 645 2405 665
rect 2425 645 2430 665
rect 2400 635 2430 645
rect 2505 655 2535 665
rect 2505 635 2510 655
rect 2530 635 2535 655
rect 2505 625 2535 635
rect 1040 565 1450 580
rect 920 525 935 550
rect 1040 525 1055 565
rect 1435 545 1450 565
rect 1790 545 1805 580
rect 1435 530 1805 545
rect 920 510 1055 525
rect 1790 420 1805 530
rect 1895 420 1910 580
rect 210 360 225 375
rect 315 360 330 375
rect 1790 305 1805 320
rect 1895 305 1910 320
<< polycont >>
rect -545 845 -525 865
rect 325 915 345 935
rect 645 915 665 935
rect -350 655 -330 675
rect 1035 850 1055 870
rect 1905 920 1925 940
rect 1230 660 1250 680
rect 2405 645 2425 665
rect 2510 635 2530 655
<< locali >>
rect -790 1215 -770 1270
rect -790 1210 -710 1215
rect -790 1140 -780 1210
rect -760 1140 -740 1210
rect -720 1140 -710 1210
rect -790 1135 -710 1140
rect -685 1210 -645 1215
rect -685 1140 -675 1210
rect -655 1140 -645 1210
rect -685 1135 -645 1140
rect -665 1085 -645 1135
rect -430 1140 -410 1210
rect -160 1140 -140 1210
rect -60 1180 130 1200
rect -60 1140 -40 1180
rect 110 1140 130 1180
rect 170 1140 190 1210
rect 790 1220 810 1275
rect 790 1215 870 1220
rect 790 1145 800 1215
rect 820 1145 840 1215
rect 860 1145 870 1215
rect 790 1140 870 1145
rect 895 1215 935 1220
rect 895 1145 905 1215
rect 925 1145 935 1215
rect 895 1140 935 1145
rect -430 1135 -350 1140
rect -665 1065 -525 1085
rect -665 1045 -645 1065
rect -790 1040 -710 1045
rect -790 970 -780 1040
rect -760 970 -740 1040
rect -720 970 -710 1040
rect -790 965 -710 970
rect -685 1040 -645 1045
rect -685 970 -675 1040
rect -655 970 -645 1040
rect -685 965 -645 970
rect -790 935 -770 965
rect -545 875 -525 1065
rect -430 1065 -420 1135
rect -400 1065 -380 1135
rect -360 1065 -350 1135
rect -430 1060 -350 1065
rect -325 1135 -245 1140
rect -325 1065 -315 1135
rect -295 1065 -275 1135
rect -255 1065 -245 1135
rect -325 1060 -245 1065
rect -220 1135 -100 1140
rect -220 1065 -210 1135
rect -190 1065 -170 1135
rect -150 1065 -130 1135
rect -110 1065 -100 1135
rect -220 1060 -100 1065
rect -80 1135 -40 1140
rect -80 1065 -70 1135
rect -50 1065 -40 1135
rect -80 1060 -40 1065
rect -15 1135 65 1140
rect -15 1065 -5 1135
rect 15 1065 35 1135
rect 55 1065 65 1135
rect -15 1060 65 1065
rect 90 1135 130 1140
rect 90 1065 100 1135
rect 120 1065 130 1135
rect 90 1060 130 1065
rect 150 1135 190 1140
rect 150 1065 160 1135
rect 180 1065 190 1135
rect 150 1060 190 1065
rect 385 1065 405 1120
rect 915 1090 935 1140
rect 1150 1145 1170 1215
rect 1420 1145 1440 1215
rect 1520 1185 1710 1205
rect 1520 1145 1540 1185
rect 1690 1145 1710 1185
rect 1750 1145 1770 1215
rect 1150 1140 1230 1145
rect 915 1070 1055 1090
rect 385 1060 465 1065
rect -295 1035 -275 1060
rect -80 1035 -60 1060
rect -295 1015 -60 1035
rect 15 935 35 1060
rect 385 990 395 1060
rect 415 990 435 1060
rect 455 990 465 1060
rect 385 985 465 990
rect 490 1060 530 1065
rect 490 990 500 1060
rect 520 990 530 1060
rect 915 1050 935 1070
rect 490 985 530 990
rect 315 935 355 945
rect -390 915 325 935
rect 345 915 355 935
rect -390 875 -370 915
rect -80 875 -60 915
rect 315 905 355 915
rect 510 935 530 985
rect 790 1045 870 1050
rect 790 975 800 1045
rect 820 975 840 1045
rect 860 975 870 1045
rect 790 970 870 975
rect 895 1045 935 1050
rect 895 975 905 1045
rect 925 975 935 1045
rect 895 970 935 975
rect 635 935 675 945
rect 510 915 645 935
rect 665 915 675 935
rect 790 940 810 970
rect 510 895 530 915
rect 635 905 675 915
rect 385 890 465 895
rect -745 805 -725 860
rect -550 865 -520 875
rect -550 845 -545 865
rect -525 845 -520 865
rect -550 835 -520 845
rect -450 870 -410 875
rect -745 800 -665 805
rect -745 730 -735 800
rect -715 730 -695 800
rect -675 730 -665 800
rect -745 725 -665 730
rect -640 800 -600 805
rect -640 730 -630 800
rect -610 730 -600 800
rect -450 800 -440 870
rect -420 800 -410 870
rect -450 795 -410 800
rect -390 870 -350 875
rect -390 800 -380 870
rect -360 800 -350 870
rect -390 795 -350 800
rect -325 870 -245 875
rect -325 800 -315 870
rect -295 800 -275 870
rect -255 800 -245 870
rect -325 795 -245 800
rect -220 870 -100 875
rect -220 800 -210 870
rect -190 800 -170 870
rect -150 800 -130 870
rect -110 800 -100 870
rect -220 795 -100 800
rect -80 870 -40 875
rect -80 800 -70 870
rect -50 800 -40 870
rect -80 795 -40 800
rect -15 870 65 875
rect -15 800 -5 870
rect 15 800 35 870
rect 55 800 65 870
rect -15 795 65 800
rect 90 870 170 875
rect 90 800 100 870
rect 120 800 140 870
rect 160 800 170 870
rect 245 845 275 855
rect 245 825 250 845
rect 270 825 275 845
rect 245 815 275 825
rect 385 820 395 890
rect 415 820 435 890
rect 455 820 465 890
rect 385 815 465 820
rect 490 890 530 895
rect 490 820 500 890
rect 520 820 530 890
rect 490 815 530 820
rect 1035 880 1055 1070
rect 1150 1070 1160 1140
rect 1180 1070 1200 1140
rect 1220 1070 1230 1140
rect 1150 1065 1230 1070
rect 1255 1140 1335 1145
rect 1255 1070 1265 1140
rect 1285 1070 1305 1140
rect 1325 1070 1335 1140
rect 1255 1065 1335 1070
rect 1360 1140 1480 1145
rect 1360 1070 1370 1140
rect 1390 1070 1410 1140
rect 1430 1070 1450 1140
rect 1470 1070 1480 1140
rect 1360 1065 1480 1070
rect 1500 1140 1540 1145
rect 1500 1070 1510 1140
rect 1530 1070 1540 1140
rect 1500 1065 1540 1070
rect 1565 1140 1645 1145
rect 1565 1070 1575 1140
rect 1595 1070 1615 1140
rect 1635 1070 1645 1140
rect 1565 1065 1645 1070
rect 1670 1140 1710 1145
rect 1670 1070 1680 1140
rect 1700 1070 1710 1140
rect 1670 1065 1710 1070
rect 1730 1140 1770 1145
rect 1730 1070 1740 1140
rect 1760 1070 1770 1140
rect 1730 1065 1770 1070
rect 1965 1070 1985 1125
rect 1965 1065 2045 1070
rect 1285 1040 1305 1065
rect 1500 1040 1520 1065
rect 1285 1020 1520 1040
rect 1595 940 1615 1065
rect 1965 995 1975 1065
rect 1995 995 2015 1065
rect 2035 995 2045 1065
rect 1965 990 2045 995
rect 2070 1065 2110 1070
rect 2070 995 2080 1065
rect 2100 995 2110 1065
rect 2070 990 2110 995
rect 1895 940 1935 950
rect 1190 920 1905 940
rect 1925 920 1935 940
rect 1190 880 1210 920
rect 1500 880 1520 920
rect 1895 910 1935 920
rect 2090 940 2110 990
rect 2320 1015 2340 1065
rect 2610 1015 2630 1065
rect 2320 1010 2400 1015
rect 2175 940 2255 960
rect 2090 920 2255 940
rect 2320 940 2330 1010
rect 2350 940 2370 1010
rect 2390 940 2400 1010
rect 2320 935 2400 940
rect 2425 1010 2505 1015
rect 2425 940 2435 1010
rect 2455 940 2475 1010
rect 2495 940 2505 1010
rect 2425 935 2505 940
rect 2530 1010 2570 1015
rect 2530 940 2540 1010
rect 2560 940 2570 1010
rect 2530 935 2570 940
rect 2590 1010 2630 1015
rect 2590 940 2600 1010
rect 2620 940 2630 1010
rect 2590 935 2630 940
rect 2090 900 2110 920
rect 2175 905 2255 920
rect 2530 900 2550 935
rect 2660 900 2775 910
rect 1965 895 2045 900
rect 90 795 170 800
rect -450 765 -430 795
rect -160 765 -140 795
rect 150 765 170 795
rect -640 725 -600 730
rect -620 675 -600 725
rect 250 715 270 815
rect 385 765 405 815
rect 835 810 855 865
rect 1030 870 1060 880
rect 1030 850 1035 870
rect 1055 850 1060 870
rect 1030 840 1060 850
rect 1130 875 1170 880
rect 835 805 915 810
rect 835 735 845 805
rect 865 735 885 805
rect 905 735 915 805
rect 835 730 915 735
rect 940 805 980 810
rect 940 735 950 805
rect 970 735 980 805
rect 1130 805 1140 875
rect 1160 805 1170 875
rect 1130 800 1170 805
rect 1190 875 1230 880
rect 1190 805 1200 875
rect 1220 805 1230 875
rect 1190 800 1230 805
rect 1255 875 1335 880
rect 1255 805 1265 875
rect 1285 805 1305 875
rect 1325 805 1335 875
rect 1255 800 1335 805
rect 1360 875 1480 880
rect 1360 805 1370 875
rect 1390 805 1410 875
rect 1430 805 1450 875
rect 1470 805 1480 875
rect 1360 800 1480 805
rect 1500 875 1540 880
rect 1500 805 1510 875
rect 1530 805 1540 875
rect 1500 800 1540 805
rect 1565 875 1645 880
rect 1565 805 1575 875
rect 1595 805 1615 875
rect 1635 805 1645 875
rect 1565 800 1645 805
rect 1670 875 1750 880
rect 1670 805 1680 875
rect 1700 805 1720 875
rect 1740 805 1750 875
rect 1825 850 1855 860
rect 1825 830 1830 850
rect 1850 830 1855 850
rect 1825 820 1855 830
rect 1965 825 1975 895
rect 1995 825 2015 895
rect 2035 825 2045 895
rect 1965 820 2045 825
rect 2070 895 2110 900
rect 2070 825 2080 895
rect 2100 825 2110 895
rect 2455 880 2775 900
rect 2455 840 2475 880
rect 2660 855 2775 880
rect 2070 820 2110 825
rect 2320 835 2400 840
rect 1670 800 1750 805
rect 1130 770 1150 800
rect 1420 770 1440 800
rect 1730 770 1750 800
rect 940 730 980 735
rect 125 695 415 715
rect -355 675 -325 685
rect -620 655 -350 675
rect -330 655 -325 675
rect -620 635 -600 655
rect -355 645 -325 655
rect 125 665 145 695
rect 395 665 415 695
rect 125 660 205 665
rect -745 630 -665 635
rect -745 560 -735 630
rect -715 560 -695 630
rect -675 560 -665 630
rect -745 555 -665 560
rect -640 630 -600 635
rect -640 560 -630 630
rect -610 560 -600 630
rect 125 590 135 660
rect 155 590 175 660
rect 195 590 205 660
rect 125 585 205 590
rect 230 660 310 665
rect 230 590 240 660
rect 260 590 280 660
rect 300 590 310 660
rect 230 585 310 590
rect 335 660 415 665
rect 335 590 345 660
rect 365 590 385 660
rect 405 590 415 660
rect 960 680 980 730
rect 1830 720 1850 820
rect 1965 770 1985 820
rect 2320 765 2330 835
rect 2350 765 2370 835
rect 2390 765 2400 835
rect 2320 760 2400 765
rect 2425 835 2505 840
rect 2425 765 2435 835
rect 2455 765 2475 835
rect 2495 765 2505 835
rect 2425 760 2505 765
rect 2530 835 2610 840
rect 2530 765 2540 835
rect 2560 765 2580 835
rect 2600 765 2610 835
rect 2530 760 2610 765
rect 1705 700 1995 720
rect 1225 680 1255 690
rect 960 660 1230 680
rect 1250 660 1255 680
rect 960 640 980 660
rect 1225 650 1255 660
rect 1705 670 1725 700
rect 1975 670 1995 700
rect 2320 715 2340 760
rect 2590 715 2610 760
rect 1705 665 1785 670
rect 335 585 415 590
rect 835 635 915 640
rect -640 555 -600 560
rect -745 515 -725 555
rect 250 525 270 585
rect 835 565 845 635
rect 865 565 885 635
rect 905 565 915 635
rect 835 560 915 565
rect 940 635 980 640
rect 940 565 950 635
rect 970 565 980 635
rect 1705 595 1715 665
rect 1735 595 1755 665
rect 1775 595 1785 665
rect 1705 590 1785 595
rect 1810 665 1890 670
rect 1810 595 1820 665
rect 1840 595 1860 665
rect 1880 595 1890 665
rect 1810 590 1890 595
rect 1915 665 1995 670
rect 2400 665 2430 675
rect 1915 595 1925 665
rect 1945 595 1965 665
rect 1985 595 1995 665
rect 1915 590 1995 595
rect 2245 645 2405 665
rect 2425 645 2430 665
rect 940 560 980 565
rect 165 505 705 525
rect 165 465 185 505
rect 105 460 145 465
rect 105 390 115 460
rect 135 390 145 460
rect 105 385 145 390
rect 165 460 205 465
rect 165 390 175 460
rect 195 390 205 460
rect 165 385 205 390
rect 230 460 310 465
rect 230 390 240 460
rect 260 390 280 460
rect 300 390 310 460
rect 230 385 310 390
rect 335 460 415 465
rect 335 390 345 460
rect 365 390 385 460
rect 405 390 415 460
rect 685 450 705 505
rect 835 520 855 560
rect 1830 530 1850 590
rect 2245 530 2265 645
rect 2400 635 2430 645
rect 2505 655 2535 665
rect 2505 635 2510 655
rect 2530 635 2535 655
rect 2505 625 2535 635
rect 1745 510 2265 530
rect 685 430 1615 450
rect 335 385 415 390
rect 105 350 125 385
rect 395 350 415 385
rect 1595 265 1615 430
rect 1745 410 1765 510
rect 1685 405 1725 410
rect 1685 335 1695 405
rect 1715 335 1725 405
rect 1685 330 1725 335
rect 1745 405 1785 410
rect 1745 335 1755 405
rect 1775 335 1785 405
rect 1745 330 1785 335
rect 1810 405 1890 410
rect 1810 335 1820 405
rect 1840 335 1860 405
rect 1880 335 1890 405
rect 1810 330 1890 335
rect 1915 405 1995 410
rect 1915 335 1925 405
rect 1945 335 1965 405
rect 1985 335 1995 405
rect 1915 330 1995 335
rect 1685 295 1705 330
rect 1975 295 1995 330
rect 2510 265 2530 625
rect 1595 245 1665 265
rect 1645 240 1665 245
rect 1725 245 1955 265
rect 1725 240 1745 245
rect 1645 220 1745 240
rect 1935 235 1955 245
rect 2015 245 2530 265
rect 2015 235 2035 245
rect 1935 215 2035 235
<< viali >>
rect -790 1270 -770 1290
rect 790 1275 810 1295
rect -430 1210 -410 1230
rect -160 1210 -140 1230
rect 170 1210 190 1230
rect -790 915 -770 935
rect -745 860 -725 880
rect 385 1120 405 1140
rect 1150 1215 1170 1235
rect 1420 1215 1440 1235
rect 1750 1215 1770 1235
rect 790 920 810 940
rect 250 825 270 845
rect 835 865 855 885
rect 1965 1125 1985 1145
rect 2320 1065 2340 1085
rect 2610 1065 2630 1085
rect -450 745 -430 765
rect -160 745 -140 765
rect 150 745 170 765
rect 385 745 405 765
rect 1830 830 1850 850
rect 1130 750 1150 770
rect 1420 750 1440 770
rect 1730 750 1750 770
rect 1965 750 1985 770
rect 2320 695 2340 715
rect 2590 695 2610 715
rect -745 495 -725 515
rect 835 500 855 520
rect 105 330 125 350
rect 395 330 415 350
rect 1685 275 1705 295
rect 1975 275 1995 295
<< metal1 >>
rect 535 1295 980 1300
rect -835 1290 -600 1295
rect -835 1270 -790 1290
rect -770 1270 -600 1290
rect -835 1265 -600 1270
rect -630 1235 -600 1265
rect 535 1275 790 1295
rect 810 1275 980 1295
rect 535 1270 980 1275
rect -630 1230 370 1235
rect -630 1210 -430 1230
rect -410 1210 -160 1230
rect -140 1210 170 1230
rect 190 1210 370 1230
rect -630 1205 370 1210
rect -835 935 -755 940
rect -835 915 -790 935
rect -770 915 -755 935
rect -835 910 -755 915
rect -835 520 -805 910
rect -630 885 -600 1205
rect -790 880 -600 885
rect -790 860 -745 880
rect -725 860 -600 880
rect -790 855 -600 860
rect 250 855 270 1205
rect 340 1145 370 1205
rect 535 1145 565 1270
rect 340 1140 565 1145
rect 340 1120 385 1140
rect 405 1120 565 1140
rect 340 1115 565 1120
rect 950 1240 980 1270
rect 950 1235 1950 1240
rect 950 1215 1150 1235
rect 1170 1215 1420 1235
rect 1440 1215 1750 1235
rect 1770 1215 1950 1235
rect 950 1210 1950 1215
rect 745 940 825 945
rect 745 920 790 940
rect 810 920 825 940
rect 745 915 825 920
rect 245 845 275 855
rect 245 825 250 845
rect 270 825 275 845
rect 245 815 275 825
rect 745 770 775 915
rect 950 890 980 1210
rect 790 885 980 890
rect 790 865 835 885
rect 855 865 980 885
rect 790 860 980 865
rect 1830 860 1850 1210
rect 1920 1150 1950 1210
rect 1920 1145 2260 1150
rect 1920 1125 1965 1145
rect 1985 1125 2260 1145
rect 1920 1120 2260 1125
rect 2230 1090 2260 1120
rect 2230 1085 2655 1090
rect 2230 1065 2320 1085
rect 2340 1065 2610 1085
rect 2630 1065 2655 1085
rect 2230 1060 2655 1065
rect 1825 850 1855 860
rect 1825 830 1830 850
rect 1850 830 1855 850
rect 1825 820 1855 830
rect -470 765 775 770
rect -470 745 -450 765
rect -430 745 -160 765
rect -140 745 150 765
rect 170 745 385 765
rect 405 745 775 765
rect -470 740 775 745
rect -470 520 -440 740
rect 745 525 775 740
rect 1110 770 2145 775
rect 1110 750 1130 770
rect 1150 750 1420 770
rect 1440 750 1730 770
rect 1750 750 1965 770
rect 1985 750 2145 770
rect 1110 745 2145 750
rect 1110 525 1140 745
rect 2305 715 2660 720
rect 2305 695 2320 715
rect 2340 695 2590 715
rect 2610 695 2660 715
rect 2305 690 2660 695
rect 2305 685 2350 690
rect 745 520 1670 525
rect -835 515 90 520
rect -835 495 -745 515
rect -725 495 90 515
rect 745 500 835 520
rect 855 500 1670 520
rect 745 495 1670 500
rect -835 490 90 495
rect 60 355 90 490
rect 60 350 430 355
rect 60 330 105 350
rect 125 330 395 350
rect 415 330 430 350
rect 60 325 430 330
rect 1640 300 1670 495
rect 2305 360 2335 685
rect 2035 330 2335 360
rect 2035 300 2065 330
rect 1640 295 2065 300
rect 1640 275 1685 295
rect 1705 275 1975 295
rect 1995 275 2065 295
rect 1640 270 2065 275
<< labels >>
flabel metal1 -820 1270 -805 1285 0 FreeSans 80 0 0 0 Vdd
port 10 nsew
flabel metal1 -830 495 -810 515 0 FreeSans 80 0 0 0 Vss
port 0 nsew
flabel poly 645 655 670 680 0 FreeSans 160 0 0 0 C
port 31 nsew
flabel poly -785 640 -760 665 0 FreeSans 160 0 0 0 B
port 33 nsew
flabel poly -830 1050 -805 1075 0 FreeSans 160 0 0 0 A
port 34 nsew
flabel locali 2200 930 2205 935 0 FreeSans 160 0 0 0 SUM
port 43 nsew
flabel locali 2710 875 2735 890 0 FreeSans 160 0 0 0 CARRY
port 46 nsew
<< end >>

magic
tech sky130A
timestamp 1766487272
<< nwell >>
rect -270 180 200 460
<< nmos >>
rect -80 0 -65 100
rect 45 0 60 100
<< pmos >>
rect -80 200 -65 400
rect 65 200 80 400
<< ndiff >>
rect -130 85 -80 100
rect -130 15 -115 85
rect -95 15 -80 85
rect -130 0 -80 15
rect -65 85 45 100
rect -65 15 -50 85
rect -30 15 10 85
rect 30 15 45 85
rect -65 0 45 15
rect 60 85 105 100
rect 60 15 75 85
rect 95 15 105 85
rect 60 0 105 15
<< pdiff >>
rect -130 385 -80 400
rect -130 215 -115 385
rect -95 215 -80 385
rect -130 200 -80 215
rect -65 385 -15 400
rect -65 215 -50 385
rect -30 215 -15 385
rect -65 200 -15 215
rect 15 385 65 400
rect 15 215 30 385
rect 50 215 65 385
rect 15 200 65 215
rect 80 385 130 400
rect 80 215 95 385
rect 120 215 130 385
rect 80 200 130 215
<< ndiffc >>
rect -115 15 -95 85
rect -50 15 -30 85
rect 10 15 30 85
rect 75 15 95 85
<< pdiffc >>
rect -115 215 -95 385
rect -50 215 -30 385
rect 30 215 50 385
rect 95 215 120 385
<< psubdiff >>
rect -185 85 -130 100
rect -185 15 -175 85
rect -155 15 -130 85
rect -185 0 -130 15
rect 105 85 145 100
rect 105 15 115 85
rect 135 15 145 85
rect 105 0 145 15
<< nsubdiff >>
rect -185 385 -130 400
rect -185 215 -175 385
rect -155 215 -130 385
rect -185 200 -130 215
rect 130 385 180 400
rect 130 215 140 385
rect 170 215 180 385
rect 130 200 180 215
<< psubdiffcont >>
rect -175 15 -155 85
rect 115 15 135 85
<< nsubdiffcont >>
rect -175 215 -155 385
rect 140 215 170 385
<< poly >>
rect -80 400 -65 460
rect 65 400 80 460
rect -80 145 -65 200
rect 65 145 80 200
rect -200 130 -65 145
rect -80 100 -65 130
rect 45 130 80 145
rect 45 100 60 130
rect -80 -15 -65 0
rect 45 -36 60 0
rect -200 -51 60 -36
<< locali >>
rect -185 390 -165 420
rect -50 390 -30 420
rect 160 390 180 420
rect -185 385 -145 390
rect -185 215 -175 385
rect -155 215 -145 385
rect -185 210 -145 215
rect -125 385 -85 390
rect -125 215 -115 385
rect -95 215 -85 385
rect -125 180 -85 215
rect -60 385 -20 390
rect -60 215 -50 385
rect -30 215 -20 385
rect -60 210 -20 215
rect 20 385 60 390
rect 20 215 30 385
rect 50 215 60 385
rect 20 210 60 215
rect 85 385 180 390
rect 85 215 95 385
rect 120 215 140 385
rect 170 215 180 385
rect 85 210 180 215
rect 20 180 40 210
rect -125 160 40 180
rect -185 85 -145 90
rect -185 15 -175 85
rect -155 15 -145 85
rect -185 10 -145 15
rect -125 85 -85 160
rect -125 15 -115 85
rect -95 15 -85 85
rect -125 10 -85 15
rect -60 85 40 90
rect -60 15 -50 85
rect -30 15 10 85
rect 30 15 40 85
rect -60 10 40 15
rect 65 85 145 90
rect 65 15 75 85
rect 95 15 115 85
rect 135 15 145 85
rect 65 10 145 15
rect -185 -70 -165 10
rect 125 -70 145 10
<< viali >>
rect -185 420 -165 440
rect -50 420 -30 440
rect 160 420 180 440
rect -185 -90 -165 -70
rect 125 -90 145 -70
<< metal1 >>
rect -200 440 200 445
rect -200 420 -185 440
rect -165 420 -50 440
rect -30 420 160 440
rect 180 420 200 440
rect -200 415 200 420
rect -200 -70 165 -65
rect -200 -90 -185 -70
rect -165 -90 125 -70
rect 145 -90 165 -70
rect -200 -95 165 -90
<< end >>
